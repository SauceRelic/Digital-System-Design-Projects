
module nios_count (
	clk_clk,
	reset_reset_n,
	pio_ssd_ext_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[15:0]	pio_ssd_ext_export;
endmodule
