
module nios_3pio (
	clk_clk,
	reset_reset_n,
	swin_pio_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	input	[3:0]	swin_pio_external_connection_export;
endmodule
