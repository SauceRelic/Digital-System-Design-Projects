	component nios_count is
		port (
			clk_clk            : in  std_logic                     := 'X'; -- clk
			reset_reset_n      : in  std_logic                     := 'X'; -- reset_n
			pio_ssd_ext_export : out std_logic_vector(15 downto 0)         -- export
		);
	end component nios_count;

	u0 : component nios_count
		port map (
			clk_clk            => CONNECTED_TO_clk_clk,            --         clk.clk
			reset_reset_n      => CONNECTED_TO_reset_reset_n,      --       reset.reset_n
			pio_ssd_ext_export => CONNECTED_TO_pio_ssd_ext_export  -- pio_ssd_ext.export
		);

